* Voltage Divider
V1 VIN 0 12
R1 VIN VOUT 10k
R2 VOUT 0 10k
.op
.dc V1 0 15 0.5
.end