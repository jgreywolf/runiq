* RL High-Pass Filter
V1 VIN 0 SIN(0 1 1k)
L1 VIN VOUT 10m
R1 VOUT 0 1k
.tran 0 5m
.ac dec 50 100 100k
.end