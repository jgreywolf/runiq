* RC Lowpass Filter
V1 IN 0 SIN(0 1 1k)
R1 IN OUT 10k
C1 OUT 0 1n
.tran 0 5m
.end