* LED Circuit with Current Limiting
V1 VCC 0 5
R1 VCC LED_ANODE 220
D1 LED_ANODE 0 2
.op
.dc V1 0 6 0.1
.end